module tb;
    

    half_adder DUT(x, y, s, c);
endmodule